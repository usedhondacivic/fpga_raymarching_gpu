// Computer_System.v

// Generated using ACDS version 23.1 991

`timescale 1 ps / 1 ps
module Computer_System (
		output wire [31:0] blue_shift_export,               //           blue_shift.export
		output wire [31:0] color_enables_export,            //        color_enables.export
		output wire [31:0] eye_x_export,                    //                eye_x.export
		output wire [31:0] eye_y_export,                    //                eye_y.export
		output wire [31:0] eye_z_export,                    //                eye_z.export
		output wire [31:0] fog_shift_export,                //            fog_shift.export
		output wire [31:0] green_shift_export,              //          green_shift.export
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //               hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                     .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                     .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                     .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                     .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                     .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                     .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                     .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                     .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                     .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                     .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                     .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                     .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                     .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,     //                     .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,     //                     .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,     //                     .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,     //                     .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,     //                     .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,     //                     .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                     .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                     .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                     .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                     .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                     .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                     .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                     .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                     .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                     .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                     .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                     .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                     .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                     .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                     .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                     .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                     .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                     .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                     .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,    //                     .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,   //                     .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,   //                     .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,    //                     .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                     .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                     .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //                     .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //                     .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //                     .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //                     .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,  //                     .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,  //                     .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,  //                     .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO41,  //                     .hps_io_gpio_inst_GPIO41
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,  //                     .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,  //                     .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,  //                     .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,  //                     .hps_io_gpio_inst_GPIO61
		output wire [31:0] lookat_1_1_export,               //           lookat_1_1.export
		output wire [31:0] lookat_1_2_export,               //           lookat_1_2.export
		output wire [31:0] lookat_1_3_export,               //           lookat_1_3.export
		output wire [31:0] lookat_2_1_export,               //           lookat_2_1.export
		output wire [31:0] lookat_2_2_export,               //           lookat_2_2.export
		output wire [31:0] lookat_2_3_export,               //           lookat_2_3.export
		output wire [31:0] lookat_3_1_export,               //           lookat_3_1.export
		output wire [31:0] lookat_3_2_export,               //           lookat_3_2.export
		output wire [31:0] lookat_3_3_export,               //           lookat_3_3.export
		output wire        m10k_pll_locked_export,          //      m10k_pll_locked.export
		output wire        m10k_pll_outclk0_clk,            //     m10k_pll_outclk0.clk
		output wire [14:0] memory_mem_a,                    //               memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                     .mem_ba
		output wire        memory_mem_ck,                   //                     .mem_ck
		output wire        memory_mem_ck_n,                 //                     .mem_ck_n
		output wire        memory_mem_cke,                  //                     .mem_cke
		output wire        memory_mem_cs_n,                 //                     .mem_cs_n
		output wire        memory_mem_ras_n,                //                     .mem_ras_n
		output wire        memory_mem_cas_n,                //                     .mem_cas_n
		output wire        memory_mem_we_n,                 //                     .mem_we_n
		output wire        memory_mem_reset_n,              //                     .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                     .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                     .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                     .mem_dqs_n
		output wire        memory_mem_odt,                  //                     .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                     .mem_dm
		input  wire        memory_oct_rzqin,                //                     .oct_rzqin
		output wire [31:0] red_shift_export,                //            red_shift.export
		output wire [31:0] repetition_pow_export,           //       repetition_pow.export
		input  wire        system_pll_ref_clk_clk,          //   system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset,      // system_pll_ref_reset.reset
		output wire        vga_pio_locked_export,           //       vga_pio_locked.export
		output wire        vga_pio_outclk0_clk              //      vga_pio_outclk0.clk
	);

	wire         system_pll_sys_clk_clk;                         // System_PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, blue_shift:clk, color_enables:clk, eye_x:clk, eye_y:clk, eye_z:clk, fog_shift:clk, green_shift:clk, lookat_1_1:clk, lookat_1_2:clk, lookat_1_3:clk, lookat_2_1:clk, lookat_2_2:clk, lookat_2_3:clk, lookat_3_1:clk, lookat_3_2:clk, lookat_3_3:clk, m10k_pll:refclk, mm_interconnect_0:System_PLL_sys_clk_clk, red_shift:clk, repetition_pow:clk, rst_controller:clk, rst_controller_003:clk, vga_pio:refclk]
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;           // ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awburst
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;             // ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlen
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;             // ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	wire         arm_a9_hps_h2f_lw_axi_master_wready;            // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_rid;               // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	wire         arm_a9_hps_h2f_lw_axi_master_rready;            // ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rready
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;             // ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlen
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_wid;               // ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;           // ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arcache
	wire         arm_a9_hps_h2f_lw_axi_master_wvalid;            // ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;            // ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_araddr
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;            // ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arprot
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;            // ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awprot
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;             // ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wdata
	wire         arm_a9_hps_h2f_lw_axi_master_arvalid;           // ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;           // ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awcache
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_arid;              // ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arid
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;            // ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlock
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;            // ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlock
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;            // ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;             // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	wire         arm_a9_hps_h2f_lw_axi_master_arready;           // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;             // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	wire         arm_a9_hps_h2f_lw_axi_master_awready;           // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;           // ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arburst
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;            // ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arsize
	wire         arm_a9_hps_h2f_lw_axi_master_bready;            // ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bready
	wire         arm_a9_hps_h2f_lw_axi_master_rlast;             // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	wire         arm_a9_hps_h2f_lw_axi_master_wlast;             // ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wlast
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;             // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_awid;              // ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awid
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_bid;               // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	wire         arm_a9_hps_h2f_lw_axi_master_bvalid;            // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;            // ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awsize
	wire         arm_a9_hps_h2f_lw_axi_master_awvalid;           // ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	wire         arm_a9_hps_h2f_lw_axi_master_rvalid;            // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	wire         mm_interconnect_0_lookat_1_1_s1_chipselect;     // mm_interconnect_0:lookat_1_1_s1_chipselect -> lookat_1_1:chipselect
	wire  [31:0] mm_interconnect_0_lookat_1_1_s1_readdata;       // lookat_1_1:readdata -> mm_interconnect_0:lookat_1_1_s1_readdata
	wire   [1:0] mm_interconnect_0_lookat_1_1_s1_address;        // mm_interconnect_0:lookat_1_1_s1_address -> lookat_1_1:address
	wire         mm_interconnect_0_lookat_1_1_s1_write;          // mm_interconnect_0:lookat_1_1_s1_write -> lookat_1_1:write_n
	wire  [31:0] mm_interconnect_0_lookat_1_1_s1_writedata;      // mm_interconnect_0:lookat_1_1_s1_writedata -> lookat_1_1:writedata
	wire         mm_interconnect_0_lookat_1_2_s1_chipselect;     // mm_interconnect_0:lookat_1_2_s1_chipselect -> lookat_1_2:chipselect
	wire  [31:0] mm_interconnect_0_lookat_1_2_s1_readdata;       // lookat_1_2:readdata -> mm_interconnect_0:lookat_1_2_s1_readdata
	wire   [1:0] mm_interconnect_0_lookat_1_2_s1_address;        // mm_interconnect_0:lookat_1_2_s1_address -> lookat_1_2:address
	wire         mm_interconnect_0_lookat_1_2_s1_write;          // mm_interconnect_0:lookat_1_2_s1_write -> lookat_1_2:write_n
	wire  [31:0] mm_interconnect_0_lookat_1_2_s1_writedata;      // mm_interconnect_0:lookat_1_2_s1_writedata -> lookat_1_2:writedata
	wire         mm_interconnect_0_lookat_1_3_s1_chipselect;     // mm_interconnect_0:lookat_1_3_s1_chipselect -> lookat_1_3:chipselect
	wire  [31:0] mm_interconnect_0_lookat_1_3_s1_readdata;       // lookat_1_3:readdata -> mm_interconnect_0:lookat_1_3_s1_readdata
	wire   [1:0] mm_interconnect_0_lookat_1_3_s1_address;        // mm_interconnect_0:lookat_1_3_s1_address -> lookat_1_3:address
	wire         mm_interconnect_0_lookat_1_3_s1_write;          // mm_interconnect_0:lookat_1_3_s1_write -> lookat_1_3:write_n
	wire  [31:0] mm_interconnect_0_lookat_1_3_s1_writedata;      // mm_interconnect_0:lookat_1_3_s1_writedata -> lookat_1_3:writedata
	wire         mm_interconnect_0_lookat_2_3_s1_chipselect;     // mm_interconnect_0:lookat_2_3_s1_chipselect -> lookat_2_3:chipselect
	wire  [31:0] mm_interconnect_0_lookat_2_3_s1_readdata;       // lookat_2_3:readdata -> mm_interconnect_0:lookat_2_3_s1_readdata
	wire   [1:0] mm_interconnect_0_lookat_2_3_s1_address;        // mm_interconnect_0:lookat_2_3_s1_address -> lookat_2_3:address
	wire         mm_interconnect_0_lookat_2_3_s1_write;          // mm_interconnect_0:lookat_2_3_s1_write -> lookat_2_3:write_n
	wire  [31:0] mm_interconnect_0_lookat_2_3_s1_writedata;      // mm_interconnect_0:lookat_2_3_s1_writedata -> lookat_2_3:writedata
	wire         mm_interconnect_0_lookat_2_2_s1_chipselect;     // mm_interconnect_0:lookat_2_2_s1_chipselect -> lookat_2_2:chipselect
	wire  [31:0] mm_interconnect_0_lookat_2_2_s1_readdata;       // lookat_2_2:readdata -> mm_interconnect_0:lookat_2_2_s1_readdata
	wire   [1:0] mm_interconnect_0_lookat_2_2_s1_address;        // mm_interconnect_0:lookat_2_2_s1_address -> lookat_2_2:address
	wire         mm_interconnect_0_lookat_2_2_s1_write;          // mm_interconnect_0:lookat_2_2_s1_write -> lookat_2_2:write_n
	wire  [31:0] mm_interconnect_0_lookat_2_2_s1_writedata;      // mm_interconnect_0:lookat_2_2_s1_writedata -> lookat_2_2:writedata
	wire         mm_interconnect_0_lookat_2_1_s1_chipselect;     // mm_interconnect_0:lookat_2_1_s1_chipselect -> lookat_2_1:chipselect
	wire  [31:0] mm_interconnect_0_lookat_2_1_s1_readdata;       // lookat_2_1:readdata -> mm_interconnect_0:lookat_2_1_s1_readdata
	wire   [1:0] mm_interconnect_0_lookat_2_1_s1_address;        // mm_interconnect_0:lookat_2_1_s1_address -> lookat_2_1:address
	wire         mm_interconnect_0_lookat_2_1_s1_write;          // mm_interconnect_0:lookat_2_1_s1_write -> lookat_2_1:write_n
	wire  [31:0] mm_interconnect_0_lookat_2_1_s1_writedata;      // mm_interconnect_0:lookat_2_1_s1_writedata -> lookat_2_1:writedata
	wire         mm_interconnect_0_lookat_3_1_s1_chipselect;     // mm_interconnect_0:lookat_3_1_s1_chipselect -> lookat_3_1:chipselect
	wire  [31:0] mm_interconnect_0_lookat_3_1_s1_readdata;       // lookat_3_1:readdata -> mm_interconnect_0:lookat_3_1_s1_readdata
	wire   [1:0] mm_interconnect_0_lookat_3_1_s1_address;        // mm_interconnect_0:lookat_3_1_s1_address -> lookat_3_1:address
	wire         mm_interconnect_0_lookat_3_1_s1_write;          // mm_interconnect_0:lookat_3_1_s1_write -> lookat_3_1:write_n
	wire  [31:0] mm_interconnect_0_lookat_3_1_s1_writedata;      // mm_interconnect_0:lookat_3_1_s1_writedata -> lookat_3_1:writedata
	wire         mm_interconnect_0_lookat_3_3_s1_chipselect;     // mm_interconnect_0:lookat_3_3_s1_chipselect -> lookat_3_3:chipselect
	wire  [31:0] mm_interconnect_0_lookat_3_3_s1_readdata;       // lookat_3_3:readdata -> mm_interconnect_0:lookat_3_3_s1_readdata
	wire   [1:0] mm_interconnect_0_lookat_3_3_s1_address;        // mm_interconnect_0:lookat_3_3_s1_address -> lookat_3_3:address
	wire         mm_interconnect_0_lookat_3_3_s1_write;          // mm_interconnect_0:lookat_3_3_s1_write -> lookat_3_3:write_n
	wire  [31:0] mm_interconnect_0_lookat_3_3_s1_writedata;      // mm_interconnect_0:lookat_3_3_s1_writedata -> lookat_3_3:writedata
	wire         mm_interconnect_0_lookat_3_2_s1_chipselect;     // mm_interconnect_0:lookat_3_2_s1_chipselect -> lookat_3_2:chipselect
	wire  [31:0] mm_interconnect_0_lookat_3_2_s1_readdata;       // lookat_3_2:readdata -> mm_interconnect_0:lookat_3_2_s1_readdata
	wire   [1:0] mm_interconnect_0_lookat_3_2_s1_address;        // mm_interconnect_0:lookat_3_2_s1_address -> lookat_3_2:address
	wire         mm_interconnect_0_lookat_3_2_s1_write;          // mm_interconnect_0:lookat_3_2_s1_write -> lookat_3_2:write_n
	wire  [31:0] mm_interconnect_0_lookat_3_2_s1_writedata;      // mm_interconnect_0:lookat_3_2_s1_writedata -> lookat_3_2:writedata
	wire         mm_interconnect_0_eye_x_s1_chipselect;          // mm_interconnect_0:eye_x_s1_chipselect -> eye_x:chipselect
	wire  [31:0] mm_interconnect_0_eye_x_s1_readdata;            // eye_x:readdata -> mm_interconnect_0:eye_x_s1_readdata
	wire   [1:0] mm_interconnect_0_eye_x_s1_address;             // mm_interconnect_0:eye_x_s1_address -> eye_x:address
	wire         mm_interconnect_0_eye_x_s1_write;               // mm_interconnect_0:eye_x_s1_write -> eye_x:write_n
	wire  [31:0] mm_interconnect_0_eye_x_s1_writedata;           // mm_interconnect_0:eye_x_s1_writedata -> eye_x:writedata
	wire         mm_interconnect_0_eye_y_s1_chipselect;          // mm_interconnect_0:eye_y_s1_chipselect -> eye_y:chipselect
	wire  [31:0] mm_interconnect_0_eye_y_s1_readdata;            // eye_y:readdata -> mm_interconnect_0:eye_y_s1_readdata
	wire   [1:0] mm_interconnect_0_eye_y_s1_address;             // mm_interconnect_0:eye_y_s1_address -> eye_y:address
	wire         mm_interconnect_0_eye_y_s1_write;               // mm_interconnect_0:eye_y_s1_write -> eye_y:write_n
	wire  [31:0] mm_interconnect_0_eye_y_s1_writedata;           // mm_interconnect_0:eye_y_s1_writedata -> eye_y:writedata
	wire         mm_interconnect_0_eye_z_s1_chipselect;          // mm_interconnect_0:eye_z_s1_chipselect -> eye_z:chipselect
	wire  [31:0] mm_interconnect_0_eye_z_s1_readdata;            // eye_z:readdata -> mm_interconnect_0:eye_z_s1_readdata
	wire   [1:0] mm_interconnect_0_eye_z_s1_address;             // mm_interconnect_0:eye_z_s1_address -> eye_z:address
	wire         mm_interconnect_0_eye_z_s1_write;               // mm_interconnect_0:eye_z_s1_write -> eye_z:write_n
	wire  [31:0] mm_interconnect_0_eye_z_s1_writedata;           // mm_interconnect_0:eye_z_s1_writedata -> eye_z:writedata
	wire         mm_interconnect_0_red_shift_s1_chipselect;      // mm_interconnect_0:red_shift_s1_chipselect -> red_shift:chipselect
	wire  [31:0] mm_interconnect_0_red_shift_s1_readdata;        // red_shift:readdata -> mm_interconnect_0:red_shift_s1_readdata
	wire   [1:0] mm_interconnect_0_red_shift_s1_address;         // mm_interconnect_0:red_shift_s1_address -> red_shift:address
	wire         mm_interconnect_0_red_shift_s1_write;           // mm_interconnect_0:red_shift_s1_write -> red_shift:write_n
	wire  [31:0] mm_interconnect_0_red_shift_s1_writedata;       // mm_interconnect_0:red_shift_s1_writedata -> red_shift:writedata
	wire         mm_interconnect_0_green_shift_s1_chipselect;    // mm_interconnect_0:green_shift_s1_chipselect -> green_shift:chipselect
	wire  [31:0] mm_interconnect_0_green_shift_s1_readdata;      // green_shift:readdata -> mm_interconnect_0:green_shift_s1_readdata
	wire   [1:0] mm_interconnect_0_green_shift_s1_address;       // mm_interconnect_0:green_shift_s1_address -> green_shift:address
	wire         mm_interconnect_0_green_shift_s1_write;         // mm_interconnect_0:green_shift_s1_write -> green_shift:write_n
	wire  [31:0] mm_interconnect_0_green_shift_s1_writedata;     // mm_interconnect_0:green_shift_s1_writedata -> green_shift:writedata
	wire         mm_interconnect_0_blue_shift_s1_chipselect;     // mm_interconnect_0:blue_shift_s1_chipselect -> blue_shift:chipselect
	wire  [31:0] mm_interconnect_0_blue_shift_s1_readdata;       // blue_shift:readdata -> mm_interconnect_0:blue_shift_s1_readdata
	wire   [1:0] mm_interconnect_0_blue_shift_s1_address;        // mm_interconnect_0:blue_shift_s1_address -> blue_shift:address
	wire         mm_interconnect_0_blue_shift_s1_write;          // mm_interconnect_0:blue_shift_s1_write -> blue_shift:write_n
	wire  [31:0] mm_interconnect_0_blue_shift_s1_writedata;      // mm_interconnect_0:blue_shift_s1_writedata -> blue_shift:writedata
	wire         mm_interconnect_0_fog_shift_s1_chipselect;      // mm_interconnect_0:fog_shift_s1_chipselect -> fog_shift:chipselect
	wire  [31:0] mm_interconnect_0_fog_shift_s1_readdata;        // fog_shift:readdata -> mm_interconnect_0:fog_shift_s1_readdata
	wire   [1:0] mm_interconnect_0_fog_shift_s1_address;         // mm_interconnect_0:fog_shift_s1_address -> fog_shift:address
	wire         mm_interconnect_0_fog_shift_s1_write;           // mm_interconnect_0:fog_shift_s1_write -> fog_shift:write_n
	wire  [31:0] mm_interconnect_0_fog_shift_s1_writedata;       // mm_interconnect_0:fog_shift_s1_writedata -> fog_shift:writedata
	wire         mm_interconnect_0_color_enables_s1_chipselect;  // mm_interconnect_0:color_enables_s1_chipselect -> color_enables:chipselect
	wire  [31:0] mm_interconnect_0_color_enables_s1_readdata;    // color_enables:readdata -> mm_interconnect_0:color_enables_s1_readdata
	wire   [1:0] mm_interconnect_0_color_enables_s1_address;     // mm_interconnect_0:color_enables_s1_address -> color_enables:address
	wire         mm_interconnect_0_color_enables_s1_write;       // mm_interconnect_0:color_enables_s1_write -> color_enables:write_n
	wire  [31:0] mm_interconnect_0_color_enables_s1_writedata;   // mm_interconnect_0:color_enables_s1_writedata -> color_enables:writedata
	wire         mm_interconnect_0_repetition_pow_s1_chipselect; // mm_interconnect_0:repetition_pow_s1_chipselect -> repetition_pow:chipselect
	wire  [31:0] mm_interconnect_0_repetition_pow_s1_readdata;   // repetition_pow:readdata -> mm_interconnect_0:repetition_pow_s1_readdata
	wire   [1:0] mm_interconnect_0_repetition_pow_s1_address;    // mm_interconnect_0:repetition_pow_s1_address -> repetition_pow:address
	wire         mm_interconnect_0_repetition_pow_s1_write;      // mm_interconnect_0:repetition_pow_s1_write -> repetition_pow:write_n
	wire  [31:0] mm_interconnect_0_repetition_pow_s1_writedata;  // mm_interconnect_0:repetition_pow_s1_writedata -> repetition_pow:writedata
	wire  [31:0] arm_a9_hps_f2h_irq0_irq;                        // irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	wire  [31:0] arm_a9_hps_f2h_irq1_irq;                        // irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                 // rst_controller:reset_out -> [blue_shift:reset_n, color_enables:reset_n, eye_x:reset_n, eye_y:reset_n, eye_z:reset_n, fog_shift:reset_n, green_shift:reset_n, lookat_1_1:reset_n, lookat_1_2:reset_n, lookat_1_3:reset_n, lookat_2_1:reset_n, lookat_2_2:reset_n, lookat_2_3:reset_n, lookat_3_1:reset_n, lookat_3_2:reset_n, lookat_3_3:reset_n, mm_interconnect_0:lookat_1_1_reset_reset_bridge_in_reset_reset, red_shift:reset_n, repetition_pow:reset_n]
	wire         system_pll_reset_source_reset;                  // System_PLL:reset_source_reset -> [rst_controller:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;             // rst_controller_001:reset_out -> m10k_pll:rst
	wire         arm_a9_hps_h2f_reset_reset;                     // ARM_A9_HPS:h2f_rst_n -> [rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	wire         rst_controller_002_reset_out_reset;             // rst_controller_002:reset_out -> vga_pio:rst
	wire         rst_controller_003_reset_out_reset;             // rst_controller_003:reset_out -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	Computer_System_ARM_A9_HPS #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_a9_hps (
		.mem_a                    (memory_mem_a),                         //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                        //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                        //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                      //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                       //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                      //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                     //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                     //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                      //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                   //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                        //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                       //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                     //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                       //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                        //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                     //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),      //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),        //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),        //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),        //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),        //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),        //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),        //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),         //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),      //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),      //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),      //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),        //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),        //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),        //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),          //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),          //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),          //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),          //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),          //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),          //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),          //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),           //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),           //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),          //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),           //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),           //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),           //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),           //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),           //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),           //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),           //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),           //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),           //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),           //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),          //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),          //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),          //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),          //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),         //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),        //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),        //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),         //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),          //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),          //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),          //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),          //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),          //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),          //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),       //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),       //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),       //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_io_hps_io_gpio_inst_GPIO41),       //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),       //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),       //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),       //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),       //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (arm_a9_hps_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk              (system_pll_sys_clk_clk),               //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                     //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                     //                  .awaddr
		.h2f_AWLEN                (),                                     //                  .awlen
		.h2f_AWSIZE               (),                                     //                  .awsize
		.h2f_AWBURST              (),                                     //                  .awburst
		.h2f_AWLOCK               (),                                     //                  .awlock
		.h2f_AWCACHE              (),                                     //                  .awcache
		.h2f_AWPROT               (),                                     //                  .awprot
		.h2f_AWVALID              (),                                     //                  .awvalid
		.h2f_AWREADY              (),                                     //                  .awready
		.h2f_WID                  (),                                     //                  .wid
		.h2f_WDATA                (),                                     //                  .wdata
		.h2f_WSTRB                (),                                     //                  .wstrb
		.h2f_WLAST                (),                                     //                  .wlast
		.h2f_WVALID               (),                                     //                  .wvalid
		.h2f_WREADY               (),                                     //                  .wready
		.h2f_BID                  (),                                     //                  .bid
		.h2f_BRESP                (),                                     //                  .bresp
		.h2f_BVALID               (),                                     //                  .bvalid
		.h2f_BREADY               (),                                     //                  .bready
		.h2f_ARID                 (),                                     //                  .arid
		.h2f_ARADDR               (),                                     //                  .araddr
		.h2f_ARLEN                (),                                     //                  .arlen
		.h2f_ARSIZE               (),                                     //                  .arsize
		.h2f_ARBURST              (),                                     //                  .arburst
		.h2f_ARLOCK               (),                                     //                  .arlock
		.h2f_ARCACHE              (),                                     //                  .arcache
		.h2f_ARPROT               (),                                     //                  .arprot
		.h2f_ARVALID              (),                                     //                  .arvalid
		.h2f_ARREADY              (),                                     //                  .arready
		.h2f_RID                  (),                                     //                  .rid
		.h2f_RDATA                (),                                     //                  .rdata
		.h2f_RRESP                (),                                     //                  .rresp
		.h2f_RLAST                (),                                     //                  .rlast
		.h2f_RVALID               (),                                     //                  .rvalid
		.h2f_RREADY               (),                                     //                  .rready
		.f2h_axi_clk              (system_pll_sys_clk_clk),               //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                     //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                     //                  .awaddr
		.f2h_AWLEN                (),                                     //                  .awlen
		.f2h_AWSIZE               (),                                     //                  .awsize
		.f2h_AWBURST              (),                                     //                  .awburst
		.f2h_AWLOCK               (),                                     //                  .awlock
		.f2h_AWCACHE              (),                                     //                  .awcache
		.f2h_AWPROT               (),                                     //                  .awprot
		.f2h_AWVALID              (),                                     //                  .awvalid
		.f2h_AWREADY              (),                                     //                  .awready
		.f2h_AWUSER               (),                                     //                  .awuser
		.f2h_WID                  (),                                     //                  .wid
		.f2h_WDATA                (),                                     //                  .wdata
		.f2h_WSTRB                (),                                     //                  .wstrb
		.f2h_WLAST                (),                                     //                  .wlast
		.f2h_WVALID               (),                                     //                  .wvalid
		.f2h_WREADY               (),                                     //                  .wready
		.f2h_BID                  (),                                     //                  .bid
		.f2h_BRESP                (),                                     //                  .bresp
		.f2h_BVALID               (),                                     //                  .bvalid
		.f2h_BREADY               (),                                     //                  .bready
		.f2h_ARID                 (),                                     //                  .arid
		.f2h_ARADDR               (),                                     //                  .araddr
		.f2h_ARLEN                (),                                     //                  .arlen
		.f2h_ARSIZE               (),                                     //                  .arsize
		.f2h_ARBURST              (),                                     //                  .arburst
		.f2h_ARLOCK               (),                                     //                  .arlock
		.f2h_ARCACHE              (),                                     //                  .arcache
		.f2h_ARPROT               (),                                     //                  .arprot
		.f2h_ARVALID              (),                                     //                  .arvalid
		.f2h_ARREADY              (),                                     //                  .arready
		.f2h_ARUSER               (),                                     //                  .aruser
		.f2h_RID                  (),                                     //                  .rid
		.f2h_RDATA                (),                                     //                  .rdata
		.f2h_RRESP                (),                                     //                  .rresp
		.f2h_RLAST                (),                                     //                  .rlast
		.f2h_RVALID               (),                                     //                  .rvalid
		.f2h_RREADY               (),                                     //                  .rready
		.h2f_lw_axi_clk           (system_pll_sys_clk_clk),               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (arm_a9_hps_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (arm_a9_hps_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (arm_a9_hps_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (arm_a9_hps_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (arm_a9_hps_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (arm_a9_hps_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (arm_a9_hps_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (arm_a9_hps_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (arm_a9_hps_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (arm_a9_hps_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (arm_a9_hps_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (arm_a9_hps_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (arm_a9_hps_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (arm_a9_hps_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (arm_a9_hps_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (arm_a9_hps_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (arm_a9_hps_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (arm_a9_hps_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (arm_a9_hps_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (arm_a9_hps_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (arm_a9_hps_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (arm_a9_hps_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (arm_a9_hps_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (arm_a9_hps_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (arm_a9_hps_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (arm_a9_hps_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (arm_a9_hps_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (arm_a9_hps_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (arm_a9_hps_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (arm_a9_hps_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (arm_a9_hps_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (arm_a9_hps_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (arm_a9_hps_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (arm_a9_hps_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (arm_a9_hps_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (arm_a9_hps_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0               (arm_a9_hps_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1               (arm_a9_hps_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	Computer_System_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (),                              //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	Computer_System_blue_shift blue_shift (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_blue_shift_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_blue_shift_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_blue_shift_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_blue_shift_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_blue_shift_s1_readdata),   //                    .readdata
		.out_port   (blue_shift_export)                           // external_connection.export
	);

	Computer_System_blue_shift color_enables (
		.clk        (system_pll_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_color_enables_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_enables_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_enables_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_enables_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_enables_s1_readdata),   //                    .readdata
		.out_port   (color_enables_export)                           // external_connection.export
	);

	Computer_System_blue_shift eye_x (
		.clk        (system_pll_sys_clk_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_eye_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_eye_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_eye_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_eye_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_eye_x_s1_readdata),   //                    .readdata
		.out_port   (eye_x_export)                           // external_connection.export
	);

	Computer_System_blue_shift eye_y (
		.clk        (system_pll_sys_clk_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_eye_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_eye_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_eye_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_eye_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_eye_y_s1_readdata),   //                    .readdata
		.out_port   (eye_y_export)                           // external_connection.export
	);

	Computer_System_blue_shift eye_z (
		.clk        (system_pll_sys_clk_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_eye_z_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_eye_z_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_eye_z_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_eye_z_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_eye_z_s1_readdata),   //                    .readdata
		.out_port   (eye_z_export)                           // external_connection.export
	);

	Computer_System_blue_shift fog_shift (
		.clk        (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_fog_shift_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_fog_shift_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_fog_shift_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_fog_shift_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_fog_shift_s1_readdata),   //                    .readdata
		.out_port   (fog_shift_export)                           // external_connection.export
	);

	Computer_System_blue_shift green_shift (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_green_shift_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_green_shift_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_green_shift_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_green_shift_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_green_shift_s1_readdata),   //                    .readdata
		.out_port   (green_shift_export)                           // external_connection.export
	);

	Computer_System_blue_shift lookat_1_1 (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_lookat_1_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lookat_1_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lookat_1_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lookat_1_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lookat_1_1_s1_readdata),   //                    .readdata
		.out_port   (lookat_1_1_export)                           // external_connection.export
	);

	Computer_System_blue_shift lookat_1_2 (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_lookat_1_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lookat_1_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lookat_1_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lookat_1_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lookat_1_2_s1_readdata),   //                    .readdata
		.out_port   (lookat_1_2_export)                           // external_connection.export
	);

	Computer_System_blue_shift lookat_1_3 (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_lookat_1_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lookat_1_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lookat_1_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lookat_1_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lookat_1_3_s1_readdata),   //                    .readdata
		.out_port   (lookat_1_3_export)                           // external_connection.export
	);

	Computer_System_blue_shift lookat_2_1 (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_lookat_2_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lookat_2_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lookat_2_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lookat_2_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lookat_2_1_s1_readdata),   //                    .readdata
		.out_port   (lookat_2_1_export)                           // external_connection.export
	);

	Computer_System_blue_shift lookat_2_2 (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_lookat_2_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lookat_2_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lookat_2_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lookat_2_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lookat_2_2_s1_readdata),   //                    .readdata
		.out_port   (lookat_2_2_export)                           // external_connection.export
	);

	Computer_System_blue_shift lookat_2_3 (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_lookat_2_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lookat_2_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lookat_2_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lookat_2_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lookat_2_3_s1_readdata),   //                    .readdata
		.out_port   (lookat_2_3_export)                           // external_connection.export
	);

	Computer_System_blue_shift lookat_3_1 (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_lookat_3_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lookat_3_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lookat_3_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lookat_3_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lookat_3_1_s1_readdata),   //                    .readdata
		.out_port   (lookat_3_1_export)                           // external_connection.export
	);

	Computer_System_blue_shift lookat_3_2 (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_lookat_3_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lookat_3_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lookat_3_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lookat_3_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lookat_3_2_s1_readdata),   //                    .readdata
		.out_port   (lookat_3_2_export)                           // external_connection.export
	);

	Computer_System_blue_shift lookat_3_3 (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_lookat_3_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lookat_3_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lookat_3_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lookat_3_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lookat_3_3_s1_readdata),   //                    .readdata
		.out_port   (lookat_3_3_export)                           // external_connection.export
	);

	Computer_System_m10k_pll m10k_pll (
		.refclk   (system_pll_sys_clk_clk),             //  refclk.clk
		.rst      (rst_controller_001_reset_out_reset), //   reset.reset
		.outclk_0 (m10k_pll_outclk0_clk),               // outclk0.clk
		.locked   (m10k_pll_locked_export)              //  locked.export
	);

	Computer_System_blue_shift red_shift (
		.clk        (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_red_shift_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_red_shift_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_red_shift_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_red_shift_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_red_shift_s1_readdata),   //                    .readdata
		.out_port   (red_shift_export)                           // external_connection.export
	);

	Computer_System_blue_shift repetition_pow (
		.clk        (system_pll_sys_clk_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_repetition_pow_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_repetition_pow_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_repetition_pow_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_repetition_pow_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_repetition_pow_s1_readdata),   //                    .readdata
		.out_port   (repetition_pow_export)                           // external_connection.export
	);

	Computer_System_vga_pio vga_pio (
		.refclk   (system_pll_sys_clk_clk),             //  refclk.clk
		.rst      (rst_controller_002_reset_out_reset), //   reset.reset
		.outclk_0 (vga_pio_outclk0_clk),                // outclk0.clk
		.locked   (vga_pio_locked_export)               //  locked.export
	);

	Computer_System_mm_interconnect_0 mm_interconnect_0 (
		.ARM_A9_HPS_h2f_lw_axi_master_awid                                        (arm_a9_hps_h2f_lw_axi_master_awid),              //                                       ARM_A9_HPS_h2f_lw_axi_master.awid
		.ARM_A9_HPS_h2f_lw_axi_master_awaddr                                      (arm_a9_hps_h2f_lw_axi_master_awaddr),            //                                                                   .awaddr
		.ARM_A9_HPS_h2f_lw_axi_master_awlen                                       (arm_a9_hps_h2f_lw_axi_master_awlen),             //                                                                   .awlen
		.ARM_A9_HPS_h2f_lw_axi_master_awsize                                      (arm_a9_hps_h2f_lw_axi_master_awsize),            //                                                                   .awsize
		.ARM_A9_HPS_h2f_lw_axi_master_awburst                                     (arm_a9_hps_h2f_lw_axi_master_awburst),           //                                                                   .awburst
		.ARM_A9_HPS_h2f_lw_axi_master_awlock                                      (arm_a9_hps_h2f_lw_axi_master_awlock),            //                                                                   .awlock
		.ARM_A9_HPS_h2f_lw_axi_master_awcache                                     (arm_a9_hps_h2f_lw_axi_master_awcache),           //                                                                   .awcache
		.ARM_A9_HPS_h2f_lw_axi_master_awprot                                      (arm_a9_hps_h2f_lw_axi_master_awprot),            //                                                                   .awprot
		.ARM_A9_HPS_h2f_lw_axi_master_awvalid                                     (arm_a9_hps_h2f_lw_axi_master_awvalid),           //                                                                   .awvalid
		.ARM_A9_HPS_h2f_lw_axi_master_awready                                     (arm_a9_hps_h2f_lw_axi_master_awready),           //                                                                   .awready
		.ARM_A9_HPS_h2f_lw_axi_master_wid                                         (arm_a9_hps_h2f_lw_axi_master_wid),               //                                                                   .wid
		.ARM_A9_HPS_h2f_lw_axi_master_wdata                                       (arm_a9_hps_h2f_lw_axi_master_wdata),             //                                                                   .wdata
		.ARM_A9_HPS_h2f_lw_axi_master_wstrb                                       (arm_a9_hps_h2f_lw_axi_master_wstrb),             //                                                                   .wstrb
		.ARM_A9_HPS_h2f_lw_axi_master_wlast                                       (arm_a9_hps_h2f_lw_axi_master_wlast),             //                                                                   .wlast
		.ARM_A9_HPS_h2f_lw_axi_master_wvalid                                      (arm_a9_hps_h2f_lw_axi_master_wvalid),            //                                                                   .wvalid
		.ARM_A9_HPS_h2f_lw_axi_master_wready                                      (arm_a9_hps_h2f_lw_axi_master_wready),            //                                                                   .wready
		.ARM_A9_HPS_h2f_lw_axi_master_bid                                         (arm_a9_hps_h2f_lw_axi_master_bid),               //                                                                   .bid
		.ARM_A9_HPS_h2f_lw_axi_master_bresp                                       (arm_a9_hps_h2f_lw_axi_master_bresp),             //                                                                   .bresp
		.ARM_A9_HPS_h2f_lw_axi_master_bvalid                                      (arm_a9_hps_h2f_lw_axi_master_bvalid),            //                                                                   .bvalid
		.ARM_A9_HPS_h2f_lw_axi_master_bready                                      (arm_a9_hps_h2f_lw_axi_master_bready),            //                                                                   .bready
		.ARM_A9_HPS_h2f_lw_axi_master_arid                                        (arm_a9_hps_h2f_lw_axi_master_arid),              //                                                                   .arid
		.ARM_A9_HPS_h2f_lw_axi_master_araddr                                      (arm_a9_hps_h2f_lw_axi_master_araddr),            //                                                                   .araddr
		.ARM_A9_HPS_h2f_lw_axi_master_arlen                                       (arm_a9_hps_h2f_lw_axi_master_arlen),             //                                                                   .arlen
		.ARM_A9_HPS_h2f_lw_axi_master_arsize                                      (arm_a9_hps_h2f_lw_axi_master_arsize),            //                                                                   .arsize
		.ARM_A9_HPS_h2f_lw_axi_master_arburst                                     (arm_a9_hps_h2f_lw_axi_master_arburst),           //                                                                   .arburst
		.ARM_A9_HPS_h2f_lw_axi_master_arlock                                      (arm_a9_hps_h2f_lw_axi_master_arlock),            //                                                                   .arlock
		.ARM_A9_HPS_h2f_lw_axi_master_arcache                                     (arm_a9_hps_h2f_lw_axi_master_arcache),           //                                                                   .arcache
		.ARM_A9_HPS_h2f_lw_axi_master_arprot                                      (arm_a9_hps_h2f_lw_axi_master_arprot),            //                                                                   .arprot
		.ARM_A9_HPS_h2f_lw_axi_master_arvalid                                     (arm_a9_hps_h2f_lw_axi_master_arvalid),           //                                                                   .arvalid
		.ARM_A9_HPS_h2f_lw_axi_master_arready                                     (arm_a9_hps_h2f_lw_axi_master_arready),           //                                                                   .arready
		.ARM_A9_HPS_h2f_lw_axi_master_rid                                         (arm_a9_hps_h2f_lw_axi_master_rid),               //                                                                   .rid
		.ARM_A9_HPS_h2f_lw_axi_master_rdata                                       (arm_a9_hps_h2f_lw_axi_master_rdata),             //                                                                   .rdata
		.ARM_A9_HPS_h2f_lw_axi_master_rresp                                       (arm_a9_hps_h2f_lw_axi_master_rresp),             //                                                                   .rresp
		.ARM_A9_HPS_h2f_lw_axi_master_rlast                                       (arm_a9_hps_h2f_lw_axi_master_rlast),             //                                                                   .rlast
		.ARM_A9_HPS_h2f_lw_axi_master_rvalid                                      (arm_a9_hps_h2f_lw_axi_master_rvalid),            //                                                                   .rvalid
		.ARM_A9_HPS_h2f_lw_axi_master_rready                                      (arm_a9_hps_h2f_lw_axi_master_rready),            //                                                                   .rready
		.System_PLL_sys_clk_clk                                                   (system_pll_sys_clk_clk),                         //                                                 System_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),             // ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.lookat_1_1_reset_reset_bridge_in_reset_reset                             (rst_controller_reset_out_reset),                 //                             lookat_1_1_reset_reset_bridge_in_reset.reset
		.blue_shift_s1_address                                                    (mm_interconnect_0_blue_shift_s1_address),        //                                                      blue_shift_s1.address
		.blue_shift_s1_write                                                      (mm_interconnect_0_blue_shift_s1_write),          //                                                                   .write
		.blue_shift_s1_readdata                                                   (mm_interconnect_0_blue_shift_s1_readdata),       //                                                                   .readdata
		.blue_shift_s1_writedata                                                  (mm_interconnect_0_blue_shift_s1_writedata),      //                                                                   .writedata
		.blue_shift_s1_chipselect                                                 (mm_interconnect_0_blue_shift_s1_chipselect),     //                                                                   .chipselect
		.color_enables_s1_address                                                 (mm_interconnect_0_color_enables_s1_address),     //                                                   color_enables_s1.address
		.color_enables_s1_write                                                   (mm_interconnect_0_color_enables_s1_write),       //                                                                   .write
		.color_enables_s1_readdata                                                (mm_interconnect_0_color_enables_s1_readdata),    //                                                                   .readdata
		.color_enables_s1_writedata                                               (mm_interconnect_0_color_enables_s1_writedata),   //                                                                   .writedata
		.color_enables_s1_chipselect                                              (mm_interconnect_0_color_enables_s1_chipselect),  //                                                                   .chipselect
		.eye_x_s1_address                                                         (mm_interconnect_0_eye_x_s1_address),             //                                                           eye_x_s1.address
		.eye_x_s1_write                                                           (mm_interconnect_0_eye_x_s1_write),               //                                                                   .write
		.eye_x_s1_readdata                                                        (mm_interconnect_0_eye_x_s1_readdata),            //                                                                   .readdata
		.eye_x_s1_writedata                                                       (mm_interconnect_0_eye_x_s1_writedata),           //                                                                   .writedata
		.eye_x_s1_chipselect                                                      (mm_interconnect_0_eye_x_s1_chipselect),          //                                                                   .chipselect
		.eye_y_s1_address                                                         (mm_interconnect_0_eye_y_s1_address),             //                                                           eye_y_s1.address
		.eye_y_s1_write                                                           (mm_interconnect_0_eye_y_s1_write),               //                                                                   .write
		.eye_y_s1_readdata                                                        (mm_interconnect_0_eye_y_s1_readdata),            //                                                                   .readdata
		.eye_y_s1_writedata                                                       (mm_interconnect_0_eye_y_s1_writedata),           //                                                                   .writedata
		.eye_y_s1_chipselect                                                      (mm_interconnect_0_eye_y_s1_chipselect),          //                                                                   .chipselect
		.eye_z_s1_address                                                         (mm_interconnect_0_eye_z_s1_address),             //                                                           eye_z_s1.address
		.eye_z_s1_write                                                           (mm_interconnect_0_eye_z_s1_write),               //                                                                   .write
		.eye_z_s1_readdata                                                        (mm_interconnect_0_eye_z_s1_readdata),            //                                                                   .readdata
		.eye_z_s1_writedata                                                       (mm_interconnect_0_eye_z_s1_writedata),           //                                                                   .writedata
		.eye_z_s1_chipselect                                                      (mm_interconnect_0_eye_z_s1_chipselect),          //                                                                   .chipselect
		.fog_shift_s1_address                                                     (mm_interconnect_0_fog_shift_s1_address),         //                                                       fog_shift_s1.address
		.fog_shift_s1_write                                                       (mm_interconnect_0_fog_shift_s1_write),           //                                                                   .write
		.fog_shift_s1_readdata                                                    (mm_interconnect_0_fog_shift_s1_readdata),        //                                                                   .readdata
		.fog_shift_s1_writedata                                                   (mm_interconnect_0_fog_shift_s1_writedata),       //                                                                   .writedata
		.fog_shift_s1_chipselect                                                  (mm_interconnect_0_fog_shift_s1_chipselect),      //                                                                   .chipselect
		.green_shift_s1_address                                                   (mm_interconnect_0_green_shift_s1_address),       //                                                     green_shift_s1.address
		.green_shift_s1_write                                                     (mm_interconnect_0_green_shift_s1_write),         //                                                                   .write
		.green_shift_s1_readdata                                                  (mm_interconnect_0_green_shift_s1_readdata),      //                                                                   .readdata
		.green_shift_s1_writedata                                                 (mm_interconnect_0_green_shift_s1_writedata),     //                                                                   .writedata
		.green_shift_s1_chipselect                                                (mm_interconnect_0_green_shift_s1_chipselect),    //                                                                   .chipselect
		.lookat_1_1_s1_address                                                    (mm_interconnect_0_lookat_1_1_s1_address),        //                                                      lookat_1_1_s1.address
		.lookat_1_1_s1_write                                                      (mm_interconnect_0_lookat_1_1_s1_write),          //                                                                   .write
		.lookat_1_1_s1_readdata                                                   (mm_interconnect_0_lookat_1_1_s1_readdata),       //                                                                   .readdata
		.lookat_1_1_s1_writedata                                                  (mm_interconnect_0_lookat_1_1_s1_writedata),      //                                                                   .writedata
		.lookat_1_1_s1_chipselect                                                 (mm_interconnect_0_lookat_1_1_s1_chipselect),     //                                                                   .chipselect
		.lookat_1_2_s1_address                                                    (mm_interconnect_0_lookat_1_2_s1_address),        //                                                      lookat_1_2_s1.address
		.lookat_1_2_s1_write                                                      (mm_interconnect_0_lookat_1_2_s1_write),          //                                                                   .write
		.lookat_1_2_s1_readdata                                                   (mm_interconnect_0_lookat_1_2_s1_readdata),       //                                                                   .readdata
		.lookat_1_2_s1_writedata                                                  (mm_interconnect_0_lookat_1_2_s1_writedata),      //                                                                   .writedata
		.lookat_1_2_s1_chipselect                                                 (mm_interconnect_0_lookat_1_2_s1_chipselect),     //                                                                   .chipselect
		.lookat_1_3_s1_address                                                    (mm_interconnect_0_lookat_1_3_s1_address),        //                                                      lookat_1_3_s1.address
		.lookat_1_3_s1_write                                                      (mm_interconnect_0_lookat_1_3_s1_write),          //                                                                   .write
		.lookat_1_3_s1_readdata                                                   (mm_interconnect_0_lookat_1_3_s1_readdata),       //                                                                   .readdata
		.lookat_1_3_s1_writedata                                                  (mm_interconnect_0_lookat_1_3_s1_writedata),      //                                                                   .writedata
		.lookat_1_3_s1_chipselect                                                 (mm_interconnect_0_lookat_1_3_s1_chipselect),     //                                                                   .chipselect
		.lookat_2_1_s1_address                                                    (mm_interconnect_0_lookat_2_1_s1_address),        //                                                      lookat_2_1_s1.address
		.lookat_2_1_s1_write                                                      (mm_interconnect_0_lookat_2_1_s1_write),          //                                                                   .write
		.lookat_2_1_s1_readdata                                                   (mm_interconnect_0_lookat_2_1_s1_readdata),       //                                                                   .readdata
		.lookat_2_1_s1_writedata                                                  (mm_interconnect_0_lookat_2_1_s1_writedata),      //                                                                   .writedata
		.lookat_2_1_s1_chipselect                                                 (mm_interconnect_0_lookat_2_1_s1_chipselect),     //                                                                   .chipselect
		.lookat_2_2_s1_address                                                    (mm_interconnect_0_lookat_2_2_s1_address),        //                                                      lookat_2_2_s1.address
		.lookat_2_2_s1_write                                                      (mm_interconnect_0_lookat_2_2_s1_write),          //                                                                   .write
		.lookat_2_2_s1_readdata                                                   (mm_interconnect_0_lookat_2_2_s1_readdata),       //                                                                   .readdata
		.lookat_2_2_s1_writedata                                                  (mm_interconnect_0_lookat_2_2_s1_writedata),      //                                                                   .writedata
		.lookat_2_2_s1_chipselect                                                 (mm_interconnect_0_lookat_2_2_s1_chipselect),     //                                                                   .chipselect
		.lookat_2_3_s1_address                                                    (mm_interconnect_0_lookat_2_3_s1_address),        //                                                      lookat_2_3_s1.address
		.lookat_2_3_s1_write                                                      (mm_interconnect_0_lookat_2_3_s1_write),          //                                                                   .write
		.lookat_2_3_s1_readdata                                                   (mm_interconnect_0_lookat_2_3_s1_readdata),       //                                                                   .readdata
		.lookat_2_3_s1_writedata                                                  (mm_interconnect_0_lookat_2_3_s1_writedata),      //                                                                   .writedata
		.lookat_2_3_s1_chipselect                                                 (mm_interconnect_0_lookat_2_3_s1_chipselect),     //                                                                   .chipselect
		.lookat_3_1_s1_address                                                    (mm_interconnect_0_lookat_3_1_s1_address),        //                                                      lookat_3_1_s1.address
		.lookat_3_1_s1_write                                                      (mm_interconnect_0_lookat_3_1_s1_write),          //                                                                   .write
		.lookat_3_1_s1_readdata                                                   (mm_interconnect_0_lookat_3_1_s1_readdata),       //                                                                   .readdata
		.lookat_3_1_s1_writedata                                                  (mm_interconnect_0_lookat_3_1_s1_writedata),      //                                                                   .writedata
		.lookat_3_1_s1_chipselect                                                 (mm_interconnect_0_lookat_3_1_s1_chipselect),     //                                                                   .chipselect
		.lookat_3_2_s1_address                                                    (mm_interconnect_0_lookat_3_2_s1_address),        //                                                      lookat_3_2_s1.address
		.lookat_3_2_s1_write                                                      (mm_interconnect_0_lookat_3_2_s1_write),          //                                                                   .write
		.lookat_3_2_s1_readdata                                                   (mm_interconnect_0_lookat_3_2_s1_readdata),       //                                                                   .readdata
		.lookat_3_2_s1_writedata                                                  (mm_interconnect_0_lookat_3_2_s1_writedata),      //                                                                   .writedata
		.lookat_3_2_s1_chipselect                                                 (mm_interconnect_0_lookat_3_2_s1_chipselect),     //                                                                   .chipselect
		.lookat_3_3_s1_address                                                    (mm_interconnect_0_lookat_3_3_s1_address),        //                                                      lookat_3_3_s1.address
		.lookat_3_3_s1_write                                                      (mm_interconnect_0_lookat_3_3_s1_write),          //                                                                   .write
		.lookat_3_3_s1_readdata                                                   (mm_interconnect_0_lookat_3_3_s1_readdata),       //                                                                   .readdata
		.lookat_3_3_s1_writedata                                                  (mm_interconnect_0_lookat_3_3_s1_writedata),      //                                                                   .writedata
		.lookat_3_3_s1_chipselect                                                 (mm_interconnect_0_lookat_3_3_s1_chipselect),     //                                                                   .chipselect
		.red_shift_s1_address                                                     (mm_interconnect_0_red_shift_s1_address),         //                                                       red_shift_s1.address
		.red_shift_s1_write                                                       (mm_interconnect_0_red_shift_s1_write),           //                                                                   .write
		.red_shift_s1_readdata                                                    (mm_interconnect_0_red_shift_s1_readdata),        //                                                                   .readdata
		.red_shift_s1_writedata                                                   (mm_interconnect_0_red_shift_s1_writedata),       //                                                                   .writedata
		.red_shift_s1_chipselect                                                  (mm_interconnect_0_red_shift_s1_chipselect),      //                                                                   .chipselect
		.repetition_pow_s1_address                                                (mm_interconnect_0_repetition_pow_s1_address),    //                                                  repetition_pow_s1.address
		.repetition_pow_s1_write                                                  (mm_interconnect_0_repetition_pow_s1_write),      //                                                                   .write
		.repetition_pow_s1_readdata                                               (mm_interconnect_0_repetition_pow_s1_readdata),   //                                                                   .readdata
		.repetition_pow_s1_writedata                                              (mm_interconnect_0_repetition_pow_s1_writedata),  //                                                                   .writedata
		.repetition_pow_s1_chipselect                                             (mm_interconnect_0_repetition_pow_s1_chipselect)  //                                                                   .chipselect
	);

	Computer_System_irq_mapper irq_mapper (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq0_irq)  //    sender.irq
	);

	Computer_System_irq_mapper irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (system_pll_reset_source_reset),  // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
